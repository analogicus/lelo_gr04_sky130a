*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_GR04_BG_lpe.spi
#else
.include ../../../work/xsch/LELO_GR04_BG.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0

* From LELO_TEMP: on from the start
VDD  VDD_1V8  0 dc {AVDD}
VPWR PWRUP_1V8 0 dc {AVDD}
VPWRN PWRUP_N_1V8 0 dc 0
V0 IBP_1F7U<0> 0 dc 0.2
V1 IBP_1F7U<1> 0 dc 0.5
V2 IBP_1F7U<2> 0 dc 0.8
V3 IBP_1F7U<3> 0 dc 1.1
VLP LPI LPO dc 0

* Save temperature: temp-sweep doesn't work for some reason
BT1 vtemp 0 V=TEMPER

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
#ifdef Debug
.save all
.option savecurrents=all
#endif

.save v(LPI)
.save i(VDD)
.save v(xdut.VX)
.save v(xdut.VY)
.save v(xdut.VD2)

* Save current probes
.save i(V0)
.save i(V1)
.save i(V2)
.save i(V3)

* Save temp
.save v(VTEMP)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 5n 5u 0
op

* -45 is gold standard
dc TEMP -55 125 5
write
quit


.endc

.end
